module function5(A0,A1,B0,f);
    input A0,A1,B0;
    output f;
    assign f = (A0&B0)|A1;
endmodule
